module fulladd(
        input a,
        input b,
        input c,
        output reg sum,
        output reg carry
    );
    always @ (*) begin
        sum=a^b^c;
        carry= (a&b) | c&(a^b);
    end
endmodule

module cla(
    input [3:0] a,b,
    input cin,
    output [3:0] sum,
    output cout
    );
    wire [3:0] p,c,g;
    assign p = a^b;
    assign g= a&b;
    
    assign c[0]=cin;
    assign c[1]= g[0] | (p[0]&c[0]);
    assign c[2]=g[1] | (p[1]&g[0]) | (p[1]&p[0]&c[0]);
    assign c[3]= g[2] | (p[2]&g[1]) |(p[2]&p[1]&g[0])| (p[2]&p[1]&p[0]&c[0]);
    assign cout=g[3] | (p[3]&g[2]) | (p[3]&p[2]&g[1]) |(p[3]&p[2]&p[1]&g[0])| (p[3]&p[2]&p[1]&p[0]&c[0]);
    assign sum= p^c;
endmodule
